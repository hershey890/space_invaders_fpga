`include "parameter_def.v"

module top_module (

);

//controls->state->state_to_display->display

endmodule