/*
 *  block_clk - clocks speed at which blocks move lower
 *      if there is time, gradually speed this up
 *  laser_clk - speed at which lasers move
 *  player_move_clk - speed at which player can move left or right
 */

module top_clock(
    input clk,
    input rst,
    output block_clk,
    output laser_clk,
    output player_move_clk,
);

endmodule