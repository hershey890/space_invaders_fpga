/*
 *  Takes switch inputs and routes them to state.v
 */

module controls (
    input rst,
    input[7:0] sw, //switch inputs
    input clk,
    output btn_adj,
    output btn_left_right,
    output btn_shoot,
);

endmodule